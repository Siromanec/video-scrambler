`timescale 1ps / 1ps
/*
modelsim wave
sim:/sequence_generator_switch_tb/generator_sequence_sig sim:/sequence_generator_switch_tb/enable_generator_sig sim:/sequence_generator_switch_tb/load_generator_sig sim:/sequence_generator_switch_tb/generator_sequence_out_sig sim:/sequence_generator_switch_tb/sequence_generator_inst/data_sig sim:/sequence_generator_switch_tb/sequence_generator_inst/shiftout_sig sim:/sequence_generator_switch_tb/clk_sig sim:/sequence_generator_switch_tb/reset_n_sig sim:/sequence_generator_switch_tb/bt656_sig sim:/sequence_generator_switch_tb/bt656_scramled sim:/sequence_generator_switch_tb/H_sig sim:/sequence_generator_switch_tb/V_out_sig sim:/sequence_generator_switch_tb/V_sig sim:/sequence_generator_switch_tb/cut_position sim:/sequence_generator_switch_tb/data_valid sim:/sequence_generator_switch_tb/prev_H sim:/sequence_generator_switch_tb/i sim:/sequence_generator_switch_tb/j sim:/sequence_generator_switch_tb/seed sim:/sequence_generator_switch_tb/H_rise
*/
module sequence_generator_switch_tb;

   localparam VIDEO_FILE_LOCATION = "video_f60.bin";
   //      localparam SCRAMBLED_VIDEO_FILE_LOCATION = "video_f60_scrambled.bin";
   localparam LINE_SIZE = 2 * 858;

   localparam LINE_COUNT = 525;
   //   localparam TOTAL_FRAMES = 60;
   localparam TOTAL_FRAMES = 10;
   localparam TOTAL_LINES = LINE_COUNT * TOTAL_FRAMES;
   localparam TOTAL_BYTES = LINE_SIZE * TOTAL_LINES;

   reg [31:0] generator_sequence_sig;
   wire enable_generator_sig;
   wire load_generator_sig;
   wire [9:0] generator_sequence_out_sig;



   reg clk_sig;
   reg reset_n_sig;
   reg [9:0] bt656_sig;
   wire [9:0] bt656_scramled;
   wire H_sig;
   wire V_sig;
   wire F_sig;
   reg [7:0] cut_position;
   wire data_valid;
   wire V_out_sig;

   //   wire [7:0] identifier_const_id;
   //   reg [9:0] detector_sequence_in_sig;
   //   wire [31:0] detector_sequence_out_sig;
   //   wire ready_sig;
   //   reg enable_detector;
   sequence_generator sequence_generator_inst (
      .clock(clk_sig),  // input  clock_sig
      .reseed_count(generator_sequence_sig),  // input [31:0] sequence_sig
      .enable(enable_generator_sig),  // input  enable_sig
      .load(load_generator_sig),  // input  load_sig
      .sequence_out(generator_sequence_out_sig)  // output [9:0] sequence_out_sig
   );
   // Generated by Quartus Prime Version 23.1 (Build Build 993 05/14/2024)
   // Created on Thu Apr 10 19:26:15 2025

   sequence_generator_switch sequence_generator_switch_inst (
      .clk(clk_sig),  // input  clk_sig
      .reset_n(reset_n_sig),  // input  reset_n_sig
      .H(H_sig),  // input  H_sig
      .V(V_sig),  // input  V_sig
      .bt656_stream_in(bt656_sig),  // input [9:0] bt656_stream_in_sig
      .sequence_in(generator_sequence_out_sig),  // input [9:0] sequence_in_sig
      .bt656_stream_out(bt656_scramled),  // output [9:0] bt656_stream_out_sig
      .V_out(V_out_sig),  // output  V_out_sig
      .enable_generator(enable_generator_sig),  // output  enable_generator_sig
      .load_generator(load_generator_sig)  // output  load_generator_sig
   );



   sync_parser sync_parser_inst (
      .clk(clk_sig),
      .reset_n(reset_n_sig),
      .bt656(bt656_sig),
      .H(H_sig),
      .V(V_sig),
      .F(F_sig)
   );

   //      line_rotator line_rotator_inst
   //      (
   //      	.clk(clk_sig) ,	// input  clk_sig
   //      	.reset_n(reset_n_sig) ,	// input  reset_n_sig
   //      	.data_in(bt656_sig) ,	// input [9:0] data_in_sig
   //      	.raw_cut_position(cut_position) ,	// input [7:0] raw_cut_position_sig
   //      	.V(V_sig) ,	// input  V_sig
   //      	.H(H_sig) ,	// input  H_sig
   //      	.data_out(bt656_scramled), 	// output [9:0] data_out_sig
   //      	.data_valid(data_valid)
   //      );


   //   reg [7:0] video_data [0:TOTAL_LINES-1];
   reg [7:0] video_value;
   integer fd;
   integer fd_out;

   reg prev_H;
   time i;
   time j;
   reg [31:0] seed;
   wire H_rise;
   assign H_rise = !prev_H & H_sig;

   reg [7:0] line_store[0:(LINE_SIZE - 1)];
   reg [7:0] line_store_out[0:(LINE_SIZE - 1)];
   initial begin
      //      cut_position = $random(seed) % 256;
      seed = 42;
      fd   = $fopen(VIDEO_FILE_LOCATION, "rb");
      if (fd == 0) begin
         $display("Error: Could not open file %s", VIDEO_FILE_LOCATION);
         $display("fd = %d", fd);
         $finish;
      end

      //         fd_out = $fopen(SCRAMBLED_VIDEO_FILE_LOCATION, "wb");
      //         if (fd_out == 0) begin
      //            $display("Error: Could not open file %s", SCRAMBLED_VIDEO_FILE_LOCATION);
      //            $display("fd_out = %d", fd_out);
      //            $finish;
      //         end
      cut_position = {$random(seed)} % 256;
      clk_sig = 0;
      reset_n_sig = 0;
      bt656_sig = 0;
      generator_sequence_sig = 0;
      #1;
      clk_sig = 0;
      #1;
      clk_sig = 1;
      reset_n_sig = 1;



      for (i = 0; i < TOTAL_BYTES / LINE_SIZE; i = i + 1) begin
         for (j = 0; j < LINE_SIZE; j = j + 1) begin
            $fgets(video_value, fd);
            line_store[j] = video_value;
            //            line_store_out[j] = 0;
         end

         generator_sequence_sig = generator_sequence_sig + 1;

         for (j = 0; j < LINE_SIZE; j = j + 1) begin
            if (H_rise && !V_sig) cut_position = {$random(seed)} % 256;


            //            $display("cut_position: %d", cut_position);
            video_value = line_store[j];

            bt656_sig  = {video_value, 2'b00};

            #1;
            clk_sig = 0;
            #1;
            clk_sig = 1;
            if (data_valid) line_store_out[j] = bt656_scramled[9:2];
            prev_H <= H_sig;
         end
         //            for (j= 0; j < LINE_SIZE; j = j + 1) begin
         //               video_value = line_store_out[j];
         //
         //               $fwrite(fd_out, "%c", video_value);
         //
         //            end

      end
      $fclose(fd);
      //         $fclose(fd_out);
      $stop;

   end


endmodule
